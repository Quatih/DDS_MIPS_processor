--------------------------------------------------------------
-- 
-- File             : test_environment.vhd
--
-- Related File(s)  : 
--
-- Author           : E. Molenkamp
-- Email            : e.molenkamp@utwente.nl
-- 
-- Project          : Digital system design
-- Creation Date    : August 23, 2012
-- 
-- Contents         : test environment for alu
--
-- Change Log 
--   Author         : 
--   Email          : 
--   Date           :  
--   Changes        :
--

library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
entity test_environment is
  generic (bw : natural := 5);
end test_environment;

